
module cordic20200720 (
	clk,
	areset,
	x,
	y,
	q);	

	input		clk;
	input		areset;
	input	[11:0]	x;
	input	[11:0]	y;
	output	[11:0]	q;
endmodule
